`timescale 1ns / 1ps
module top_efect4(input efect4 );
	 reg temp4;
always @(efect4) begin
		if (efect4)  temp4<= 1'b1;
	end


endmodule
