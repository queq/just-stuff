`timescale 1ns / 1ps
module top_efect1(input efect1 );
	 reg temp1;
always @(efect1) begin
		if (efect1)  temp1<= 1'b1;
	end


endmodule
