`timescale 1ns / 1ps
module top_efect2(input efect2 );
	 reg temp2;
always @(efect2) begin
		if (efect2)  temp2<= 1'b1;
	end


endmodule
