`timescale 1ns / 1ps
module top_efect5(input efect5 );
	 reg temp5;
always @(efect5) begin
		if (efect5)  temp5<= 1'b1;
	end


endmodule
